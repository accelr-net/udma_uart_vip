package model_pkg;
    `include "spi_master_bfm.sv"
endpackage